----------------------------------------------------------------------------------
-- Company:
-- Author:
-- 
-- Create Date:    
-- Design Name: 
-- Module Name:    
-- Project Name: 
-- Target Devices: 
-- Tool versions:
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
--Module Description

-- LUT for inverse((A.A')

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

library WORK ;
use work.ATISpackage.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;


entity a_inverse_lut_rom is
port(
	rst				: in std_logic ;
	clk				: in std_logic ;
	
	address_rdy		: in std_logic ;
	address			: in std_logic_Vector(7 downto 0);
	
	data_out_valid		: out std_logic ;
	data_out				: out AtA_inv_type
	);
end entity ;


architecture rtl of a_inverse_lut_rom is

signal data				: AtA_inv_type;
signal data_valid		: STD_LOGIC;

type mem is array (0 to  129) of std_logic_vector(127 downto 0);

-- the entries are scale by *2048
constant a_inverse_lut : mem :=(
						0	=> 	x"00000_155_000_000_000_155_000_000_000_0E3",
						1 	=> 	x"00000_1BB_066_FBB_066_1BB_FBB_FBB_FBB_111",
						2 	=> 	x"00000_1A4_000_FCB_000_155_000_FCB_000_106",
						3 	=> 	x"00000_1BB_F99_FBB_F99_1BB_044_FBB_044_111",
						4 	=> 	x"00000_155_000_000_000_1A4_FCB_000_FCB_106",
						5 	=> 	x"00000_155_000_000_000_155_000_000_000_100",
						6 	=> 	x"00000_155_000_000_000_1A4_034_000_034_106",
						7 	=> 	x"00000_1BB_F99_044_F99_1BB_FBB_044_FBB_111",
						8 	=> 	x"00000_1A4_000_034_000_155_000_034_000_106",
						9 	=> 	x"00000_1BB_066_044_066_1BB_044_044_044_111",
						10	=> 	x"00000_297_0AF_F29_0AF_1D4_F8A_F29_F8A_172",
						11	=> 	x"00000_255_000_F55_000_200_000_F55_000_155",
						12	=> 	x"00000_1D4_0AF_F8A_0AF_297_F29_F8A_F29_172",
						13	=> 	x"00000_1BE_069_FB1_069_1BE_FB1_FB1_FB1_13B",
						14	=> 	x"00000_1BC_06F_FC0_06F_21B_FF0_FC0_FF0_12D",
						15	=> 	x"00000_200_000_000_000_255_F55_000_F55_155",
						16	=> 	x"00000_21B_06F_FF0_06F_1BC_FC0_FF0_FC0_12D",
						17	=> 	x"00000_2AA_155_000_155_2AA_000_000_000_124",
						18	=> 	x"00000_297_F50_F29_F50_1D4_075_F29_075_172",
						19	=> 	x"00000_1A6_00C_FC1_00C_1A6_FC1_FC1_FC1_136",
						20	=> 	x"00000_1A5_000_FC3_000_155_000_FC3_000_12D",
						21	=> 	x"00000_1A6_FF3_FC1_FF3_1A6_03E_FC1_03E_136",
						22	=> 	x"00000_21B_F90_00F_F90_1BC_FC0_00F_FC0_12D",
						23	=> 	x"00000_200_000_000_000_155_000_000_000_124",
						24	=> 	x"00000_21B_06F_00F_06F_1BC_03F_00F_03F_12D",
						25	=> 	x"00000_1BC_F90_FC0_F90_21B_00F_FC0_00F_12D",
						26	=> 	x"00000_1BE_F96_FB1_F96_1BE_04E_FB1_04E_13B",
						27	=> 	x"00000_1D4_F50_F8A_F50_297_0D6_F8A_0D6_172",
						28	=> 	x"00000_2AA_EAA_000_EAA_2AA_000_000_000_124",
						29	=> 	x"00000_21B_F90_FF0_F90_1BC_03F_FF0_03F_12D",
						30	=> 	x"00000_200_000_000_000_255_0AA_000_0AA_155",
						31	=> 	x"00000_155_000_000_000_1A5_FC3_000_FC3_12D",
						32	=> 	x"00000_155_000_000_000_200_000_000_000_124",
						33	=> 	x"00000_1D4_F50_075_F50_297_F29_075_F29_172",
						34	=> 	x"00000_1A6_FF3_03E_FF3_1A6_FC1_03E_FC1_136",
						35	=> 	x"00000_1BC_06F_03F_06F_21B_00F_03F_00F_12D",
						36	=> 	x"00000_155_000_000_000_1A5_03C_000_03C_12D",
						37	=> 	x"00000_1BE_F96_04E_F96_1BE_FB1_04E_FB1_13B",
						38	=> 	x"00000_1A5_000_03C_000_155_000_03C_000_12D",
						39	=> 	x"00000_1BE_069_04E_069_1BE_04E_04E_04E_13B",
						40	=> 	x"00000_1BC_F90_03F_F90_21B_FF0_03F_FF0_12D",
						41	=> 	x"00000_1A6_00C_03E_00C_1A6_03E_03E_03E_136",
						42	=> 	x"00000_1D4_0AF_075_0AF_297_0D6_075_0D6_172",
						43	=> 	x"00000_297_F50_0D6_F50_1D4_F8A_0D6_F8A_172",
						44	=> 	x"00000_255_000_0AA_000_200_000_0AA_000_155",
						45	=> 	x"00000_297_0AF_0D6_0AF_1D4_075_0D6_075_172",
						46	=> 	x"00000_555_000_D55_000_200_000_D55_000_2AA",
						47	=> 	x"00000_333_199_E66_199_333_E66_E66_E66_266",
						48	=> 	x"00000_2B2_0BE_EFA_0BE_1DC_F71_EFA_F71_1C4",
						49	=> 	x"00000_298_0A6_F22_0A6_229_FC8_F22_FC8_19F",
						50	=> 	x"00000_2DB_049_F6D_049_26D_F24_F6D_F24_1B6",
						51	=> 	x"00000_322_0C1_F59_0C1_1D6_F91_F59_F91_183",
						52	=> 	x"00000_45D_22E_F45_22E_317_FA2_F45_FA2_174",
						53	=> 	x"00000_26D_049_F24_049_2DB_F6D_F24_F6D_1B6",
						54	=> 	x"00000_266_000_F33_000_200_000_F33_000_199",
						55	=> 	x"00000_26D_FB6_F24_FB6_2DB_092_F24_092_1B6",
						56	=> 	x"00000_317_F17_FA2_F17_317_FA2_FA2_FA2_174",
						57	=> 	x"00000_2D2_000_F87_000_200_000_F87_000_169",
						58	=> 	x"00000_317_0E8_FA2_0E8_317_05D_FA2_05D_174",
						59	=> 	x"00000_1DC_0BE_F71_0BE_2B2_EFA_F71_EFA_1C4",
						60	=> 	x"00000_1D6_0C1_F91_0C1_322_F59_F91_F59_183",
						61	=> 	x"00000_200_000_000_000_555_D55_000_D55_2AA",
						62	=> 	x"00000_229_0A6_FC8_0A6_298_F22_FC8_F22_19F",
						63	=> 	x"00000_317_22E_FA2_22E_45D_F45_FA2_F45_174",
						64	=> 	x"00000_1BE_06F_FB5_06F_21B_FED_FB5_FED_161",
						65	=> 	x"00000_200_000_000_000_266_F33_000_F33_199",
						66	=> 	x"00000_21B_06F_FED_06F_1BE_FB5_FED_FB5_161",
						67	=> 	x"00000_2AA_155_000_155_2AA_000_000_000_155",
						68	=> 	x"00000_200_000_000_000_2D2_F87_000_F87_169",
						69	=> 	x"00000_222_088_000_088_222_000_000_000_155",
						70	=> 	x"00000_317_22E_05D_22E_45D_0BA_05D_0BA_174",
						71	=> 	x"00000_2DB_FB6_092_FB6_26D_F24_092_F24_1B6",
						72	=> 	x"00000_317_0E8_05D_0E8_317_FA2_05D_FA2_174",
						73	=> 	x"00000_45D_22E_0BA_22E_317_05D_0BA_05D_174",
						74	=> 	x"00000_298_F59_F22_F59_229_037_F22_037_19F",
						75	=> 	x"00000_2B2_F41_EFA_F41_1DC_08E_EFA_08E_1C4",
						76	=> 	x"00000_333_E66_E66_E66_333_199_E66_199_266",
						77	=> 	x"00000_45D_DD1_F45_DD1_317_05D_F45_05D_174",
						78	=> 	x"00000_322_F3E_F59_F3E_1D6_06E_F59_06E_183",
						79	=> 	x"00000_2DB_FB6_F6D_FB6_26D_0DB_F6D_0DB_1B6",
						80	=> 	x"00000_1A8_00E_FB6_00E_1A8_FB6_FB6_FB6_16D",
						81	=> 	x"00000_1A7_000_FB9_000_200_000_FB9_000_161",
						82	=> 	x"00000_229_F59_037_F59_298_F22_037_F22_19F",
						83	=> 	x"00000_200_000_000_000_1A7_FB9_000_FB9_161",
						84	=> 	x"00000_222_088_000_088_222_000_000_000_155",
						85	=> 	x"00000_1A8_FF1_FB6_FF1_1A8_049_FB6_049_16D",
						86	=> 	x"00000_21B_F90_012_F90_1BE_FB5_012_FB5_161",
						87	=> 	x"00000_200_000_000_000_155_000_000_000_155",
						88	=> 	x"00000_21B_06F_012_06F_1BE_04A_012_04A_161",
						89	=> 	x"00000_222_F77_000_F77_222_000_000_000_155",
						90	=> 	x"00000_200_000_000_000_1A7_046_000_046_161",
						91	=> 	x"00000_229_0A6_037_0A6_298_0DD_037_0DD_19F",
						92	=> 	x"00000_322_F3E_0A6_F3E_1D6_F91_0A6_F91_183",
						93	=> 	x"00000_2D2_000_078_000_200_000_078_000_169",
						94	=> 	x"00000_322_0C1_0A6_0C1_1D6_06E_0A6_06E_183",
						95	=> 	x"00000_1BE_F90_FB5_F90_21B_012_FB5_012_161",
						96	=> 	x"00000_1D6_F3E_F91_F3E_322_0A6_F91_0A6_183",
						97	=> 	x"00000_317_DD1_05D_DD1_45D_F45_05D_F45_174",
						98	=> 	x"00000_222_F77_000_F77_222_000_000_000_155",
						99	=> 	x"00000_200_000_000_000_2D2_078_000_078_169",
						100	=> x"00000_1DC_F41_F71_F41_2B2_105_F71_105_1C4",
						101	=> x"00000_2AA_EAA_000_EAA_2AA_000_000_000_155",
						102	=> x"00000_21B_F90_FED_F90_1BE_04A_FED_04A_161",
						103	=> x"00000_200_000_000_000_266_0CC_000_0CC_199",
						104	=> x"00000_317_DD1_FA2_DD1_45D_0BA_FA2_0BA_174",
						105	=> x"00000_229_F59_FC8_F59_298_0DD_FC8_0DD_19F",
						106	=> x"00000_200_000_000_000_555_2AA_000_2AA_2AA",
						107	=> x"00000_45D_DD1_0BA_DD1_317_FA2_0BA_FA2_174",
						108	=> x"00000_317_F17_05D_F17_317_05D_05D_05D_174",
						109	=> x"00000_2DB_049_092_049_26D_0DB_092_0DB_1B6",
						110	=> x"00000_155_000_000_000_200_000_000_000_155",
						111	=> x"00000_1DC_F41_08E_F41_2B2_EFA_08E_EFA_1C4",
						112	=> x"00000_1A8_FF1_049_FF1_1A8_FB6_049_FB6_16D",
						113	=> x"00000_1BE_06F_04A_06F_21B_012_04A_012_161",
						114	=> x"00000_1D6_F3E_06E_F3E_322_F59_06E_F59_183",
						115	=> x"00000_1A7_000_046_000_200_000_046_000_161",
						116	=> x"00000_1D6_0C1_06E_0C1_322_0A6_06E_0A6_183",
						117	=> x"00000_333_E66_199_E66_333_E66_199_E66_266",
						118	=> x"00000_26D_FB6_0DB_FB6_2DB_F6D_0DB_F6D_1B6",
						119	=> x"00000_298_0A6_0DD_0A6_229_037_0DD_037_19F",
						120	=> x"00000_1BE_F90_04A_F90_21B_FED_04A_FED_161",
						121	=> x"00000_1A8_00E_049_00E_1A8_049_049_049_16D",
						122	=> x"00000_1DC_0BE_08E_0BE_2B2_105_08E_105_1C4",
						123	=> x"00000_2B2_F41_105_F41_1DC_F71_105_F71_1C4",
						124	=> x"00000_266_000_0CC_000_200_000_0CC_000_199",
						125	=> x"00000_2B2_0BE_105_0BE_1DC_08E_105_08E_1C4",
						126	=> x"00000_298_F59_0DD_F59_229_FC8_0DD_FC8_19F",
						127	=> x"00000_26D_049_0DB_049_2DB_092_0DB_092_1B6",
						128	=> x"00000_333_199_199_199_333_199_199_199_266",
						129	=> x"00000_555_000_2AA_000_200_000_2AA_000_2AA"						
						);	


begin

rom_proc: process(clk)
begin
	if rising_edge(clk) then
		--one clock cycle delay for timing synchronization
		data_out_valid <= data_valid;
		data_out <= data;
		
		if rst = '1' then
			data <= (others=> (others=> (others=> '0' )));
			data_valid <= '0' ;
		else
			data_valid <= address_rdy;
			if address_rdy = '1' then
				for y in -1 to 1 loop
					for x in y to 1 loop
						data(y)(x) <= a_inverse_lut(to_integer(unsigned(address)))(12*((-x+1)+(-y+1)*3+1)-1 downto 12*((-x+1)+(-y+1)*3));
					end loop;
					for x in -1 to (y-1) loop --exploiting symmetry, line is same as above, but with x-y swapped
						data(y)(x) <= a_inverse_lut(to_integer(unsigned(address)))(12*((-y+1)+(-x+1)*3+1)-1 downto 12*((-y+1)+(-x+1)*3));
					end loop;
				end loop;
				
			end if ;
		end if ;
	end if;
end process;		

end rtl;

